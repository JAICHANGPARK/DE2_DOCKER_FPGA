Library ieee;
USE ieee.std_logic_1164.ALL;

entity my_traffic_light is
	port (clk, vehicle : in std_logic;
		  led : out std_logic_vector(2 downto 0); 
		  led_side : out std_logic_vector(2 downto 0); 
		  btn : in STD_LOGIC_VECTOR(3 downto 3); 
		  ld : out STD_LOGIC_VECTOR(7 downto 2);
		  main, side : out natural range 0 to 7);
end my_traffic_light;

architecture behavior of my_traffic_light is
type statestype is (firststate, secondstate, thirdstate, fourthstate);
signal state, nextstate : statestype := firststate;
signal longtime, shorttime, long, short, timetrig, Fout : std_logic;
signal Setcount : integer;
signal S : std_logic_vector(0 to 1);
signal clr, clk3: STD_LOGIC; 


component timer is
	port (enable, clock : in std_logic;
		  SetCount : in integer;
		  Qout : buffer std_logic);
end component;

component frequency_divider is
	port (clock : in std_logic;
		  Fout : inout std_logic);
end component;

component lightsequence is
	port (VS, TL, CLK, TS : in std_logic;
		  S : buffer std_logic_vector(0 to 1)
		 );
end component;

component clkdiv is
 port(
 mclk : in STD_LOGIC;
 clr : in STD_LOGIC;
 clk190 : out STD_LOGIC;
 clk3 : out STD_LOGIC
 );
end component; 

begin

clr <= btn(3); 

U1: clkdiv
 port map (
 mclk=>clk,
 clr=>clr,
 clk3=>clk3
); 
 
--FR : frequency_divider port map (clock => clk , Fout => Fout);

Readstate:process(S)
begin
	case S is
		when "00" => state <= firststate;
		when "01" => state <= secondstate;
		when "10" => state <= thirdstate;
		when "11" => state <= fourthstate;
		when others => state <= firststate;
	end case;
end process Readstate;

StateDiag:process(state, clk)
begin
	case state is
		when firststate => 
			main <= 2#001#;
			side <= 2#100#;
			Setcount <= 16#19BFC#;
			led  <= "001";
			led_side <= "100";
			long <= '1';
			short <= '0';
		when secondstate => 
			main <= 2#010#;
			side <= 2#100#;
			Setcount <= 16#A0EE7#;
			led  <= "010";
			led_side <= "100";
			long <= '0';
			short <= '1';
		when thirdstate => 
			main <= 2#100#;
			side <= 2#001#;
			Setcount <= 16#19BFC#;
			led  <= "100";
			led_side <= "001";
			long <= '1';
			short <= '0';
		when fourthstate => 
			main <= 2#100#;
			side <= 2#010#;
			Setcount <= 16#A0EE7#;
			led  <= "100";
			led_side <= "010";
			long <= '0';
			short <= '1';
	end case;
end process;
end behavior;
